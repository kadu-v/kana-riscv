module riscv_alu (
    ports
);

endmodule
