/*---------------------------------------------------
Instructions
-----------------------------------------------------*/
/* R type--------------------------------------------*/
// add
`define INST_ADD 32'b0000000_00000_00000_000_00000_0110011
`define INST_ADD_MASK 32'b1111111_00000_00000_111_00000_1111111


/* I type--------------------------------------------*/
// addi
// `define INST_ADDI 
